library verilog;
use verilog.vl_types.all;
entity Branch_unit_vlg_check_tst is
    port(
        NextPCSrc       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Branch_unit_vlg_check_tst;
