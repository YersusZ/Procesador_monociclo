library verilog;
use verilog.vl_types.all;
entity Register_unit_vlg_vec_tst is
end Register_unit_vlg_vec_tst;
