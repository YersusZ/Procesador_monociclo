library verilog;
use verilog.vl_types.all;
entity Data_memory_vlg_vec_tst is
end Data_memory_vlg_vec_tst;
