library verilog;
use verilog.vl_types.all;
entity Branch_unit_vlg_vec_tst is
end Branch_unit_vlg_vec_tst;
