library verilog;
use verilog.vl_types.all;
entity Imm_unit_vlg_vec_tst is
end Imm_unit_vlg_vec_tst;
