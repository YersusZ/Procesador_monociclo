library verilog;
use verilog.vl_types.all;
entity Registro_32bits_vlg_vec_tst is
end Registro_32bits_vlg_vec_tst;
