library verilog;
use verilog.vl_types.all;
entity Procesador_monociclo is
    port(
        Clk             : in     vl_logic
    );
end Procesador_monociclo;
