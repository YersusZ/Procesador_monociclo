library verilog;
use verilog.vl_types.all;
entity Data_memory_vlg_check_tst is
    port(
        DataRd          : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end Data_memory_vlg_check_tst;
